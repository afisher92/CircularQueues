module Queues_tb();

Queues iQ (.clk(clk), .rst_n(rst_n), .newsmpl(newsmpl), .wrt_smpl(wrt_smpl), .smpl_out(smpl_out), .sequencing(sequencing));







endmodule
